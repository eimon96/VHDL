LIBRARY ieee;
USE ieee.std_logic_1164.all;


ENTITY mux_4to1_tb IS END mux_4to1_tb;


ARCHITECTURE LogicFunc_tb OF mux_4to1_tb IS
	component tbc is
port (
	clk : bit;
	x0, x1, x2, x3, s1, s0 : IN STD_LOGIC;
	f : OUT STD_LOGIC);
END COMPONENT;

	CONSTANT period : TIME := 50 ns;

	signal clk : BIT := '0';
	signal done : boolean := false;
	signal x0, x1, x2, x3, s1, s0 : STD_LOGIC := '0';
	signal f: STD_LOGIC;

begin
	u1 : tbc
	port map(
		clk => clk,
		x0 => x0,
		x1 => x1,
		x2 => x2,
		x3 => x3,
		s1 => s1,
		s0 => s0,
		f => f);
		
	clkprocess: process(done, clk)
		begin
			if (not done) then
				clk <= not clk after period / 2;
			end if;
	end process;
	
		
		f <= ( (NOT s1) AND (NOT s0) AND x0 ) OR ( (NOT s1) AND s0 AND x1 ) OR ( s1 AND (NOT s0) AND x2 ) OR ( s1 AND s0 AND x3 );
	
	
	testbench: process
		begin
			wait until (clk = '0');
			s1 <= '0';
			s0 <= '0';
			x0 <= '0';
			x1 <= '0';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '0';
			x1 <= '0';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '0';
			x1 <= '0';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '0';
			x1 <= '0';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '0';
			x1 <= '1';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '0';
			x1 <= '1';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '0';
			x1 <= '1';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '0';
			x1 <= '1';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '1';
			x1 <= '0';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '1';
			x1 <= '0';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '1';
			x1 <= '0';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '1';
			x1 <= '0';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '1';
			x1 <= '1';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '1';
			x1 <= '1';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '1';
			x1 <= '1';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '0';
			x0 <= '1';
			x1 <= '1';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '0';
			x1 <= '0';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '0';
			x1 <= '0';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '0';
			x1 <= '0';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '0';
			x1 <= '0';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '0';
			x1 <= '1';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '0';
			x1 <= '1';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '0';
			x1 <= '1';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '0';
			x1 <= '1';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '1';
			x1 <= '0';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '1';
			x1 <= '0';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '1';
			x1 <= '0';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '1';
			x1 <= '0';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '1';
			x1 <= '1';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '1';
			x1 <= '1';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '1';
			x1 <= '1';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '0';
			s0 <= '1';
			x0 <= '1';
			x1 <= '1';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '0';
			x1 <= '0';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '0';
			x1 <= '0';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '0';
			x1 <= '0';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '0';
			x1 <= '0';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '0';
			x1 <= '1';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '0';
			x1 <= '1';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '0';
			x1 <= '1';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '0';
			x1 <= '1';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '1';
			x1 <= '0';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '1';
			x1 <= '0';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '1';
			x1 <= '0';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '1';
			x1 <= '0';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '1';
			x1 <= '1';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '1';
			x1 <= '1';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '1';
			x1 <= '1';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '0';
			x0 <= '1';
			x1 <= '1';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '0';
			x1 <= '0';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '0';
			x1 <= '0';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '0';
			x1 <= '0';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '0';
			x1 <= '0';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '0';
			x1 <= '1';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '0';
			x1 <= '1';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '0';
			x1 <= '1';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '0';
			x1 <= '1';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '1';
			x1 <= '0';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '1';
			x1 <= '0';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '1';
			x1 <= '0';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '1';
			x1 <= '0';
			x2 <= '1';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '1';
			x1 <= '1';
			x2 <= '0';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '1';
			x1 <= '1';
			x2 <= '0';
			x3 <= '1';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '1';
			x1 <= '1';
			x2 <= '1';
			x3 <= '0';
			wait for period;
			s1 <= '1';
			s0 <= '1';
			x0 <= '1';
			x1 <= '1';
			x2 <= '1';
			x3 <= '1';
		    	wait for period;
			
			done <= true;
			wait;
		end process;
end LogicFunc_tb;

